`timescale 1ns / 1ps
module tb;
  
  wire o0, o1, o2, o3, o4, o5, o6, o7;     // 8 wires for 8 outputs 
  reg i0,i1,i2,i3,i4,i5,i6,i7;      // 8 regs for 8 inputs
  num N1(i0,i1,i2,i3,i4,i5,i6,i7,o0,o1,o2,o3,o4,o5,o6,o7);

initial //50 as arbitrary inter-input delay to begin with before we find threshold
  begin
    $dumpfile("wave.vcd");
    $dumpvars(0, tb, N1);
    i0 = 1'b0; i1 = 1'b0; i2 = 1'b1; i3 = 1'b0; i4 = 1'b1; i5 = 1'b0; i6 = 1'b0; i7 = 1'b0; // testing 00101000
    #50 i0 = 1'b0; i1 = 1'b1; i2 = 1'b0; i3 = 1'b0; i4 = 1'b1; i5 = 1'b0; i6 = 1'b0; i7 = 1'b0; // testing 01001000    
    #50 i0 = 1'b1; i1 = 1'b0; i2 = 1'b1; i3 = 1'b1; i4 = 1'b0; i5 = 1'b1; i6 = 1'b1; i7 = 1'b1; // testing 10110111    
    #50 i0 = 1'b1; i1 = 1'b0; i2 = 1'b0; i3 = 1'b0; i4 = 1'b0; i5 = 1'b0; i6 = 1'b1; i7 = 1'b1; // testing 10000011 
    #50 i0 = 1'b0; i1 = 1'b1; i2 = 1'b1; i3 = 1'b1; i4 = 1'b1; i5 = 1'b1; i6 = 1'b0; i7 = 1'b0; // testing 01111100    
    #50 i0 = 1'b0; i1 = 1'b0; i2 = 1'b0; i3 = 1'b1; i4 = 1'b0; i5 = 1'b1; i6 = 1'b0; i7 = 1'b0; // testing 00010100    
    #50 i0 = 1'b1; i1 = 1'b1; i2 = 1'b1; i3 = 1'b0; i4 = 1'b1; i5 = 1'b0; i6 = 1'b1; i7 = 1'b1; // testing 11101011    
    #50 i0 = 1'b0; i1 = 1'b1; i2 = 1'b1; i3 = 1'b0; i4 = 1'b0; i5 = 1'b0; i6 = 1'b0; i7 = 1'b1; // testing 01100001    
    #50 i0 = 1'b0; i1 = 1'b1; i2 = 1'b0; i3 = 1'b0; i4 = 1'b0; i5 = 1'b0; i6 = 1'b0; i7 = 1'b1; // testing 01000001    
    #50 i0 = 1'b0; i1 = 1'b1; i2 = 1'b1; i3 = 1'b1; i4 = 1'b1; i5 = 1'b0; i6 = 1'b1; i7 = 1'b0; // testing 01111010    
    #50 i0 = 1'b0; i1 = 1'b1; i2 = 1'b0; i3 = 1'b0; i4 = 1'b0; i5 = 1'b1; i6 = 1'b1; i7 = 1'b1; // testing 01000111    
    #50 i0 = 1'b0; i1 = 1'b1; i2 = 1'b1; i3 = 1'b0; i4 = 1'b1; i5 = 1'b1; i6 = 1'b0; i7 = 1'b1; // testing 01101101    
    #50 i0 = 1'b1; i1 = 1'b0; i2 = 1'b0; i3 = 1'b1; i4 = 1'b0; i5 = 1'b0; i6 = 1'b1; i7 = 1'b0; // testing 10010010    
    #50 i0 = 1'b0; i1 = 1'b0; i2 = 1'b1; i3 = 1'b1; i4 = 1'b0; i5 = 1'b0; i6 = 1'b0; i7 = 1'b0; // testing 00110000    
    #50 i0 = 1'b1; i1 = 1'b1; i2 = 1'b0; i3 = 1'b0; i4 = 1'b1; i5 = 1'b1; i6 = 1'b1; i7 = 1'b1; // testing 11001111    
    #50 i0 = 1'b0; i1 = 1'b0; i2 = 1'b1; i3 = 1'b1; i4 = 1'b1; i5 = 1'b0; i6 = 1'b1; i7 = 1'b0; // testing 00111010    
    #50 i0 = 1'b0; i1 = 1'b1; i2 = 1'b1; i3 = 1'b1; i4 = 1'b1; i5 = 1'b0; i6 = 1'b1; i7 = 1'b1; // testing 01111011    
    #50 i0 = 1'b1; i1 = 1'b0; i2 = 1'b0; i3 = 1'b0; i4 = 1'b0; i5 = 1'b1; i6 = 1'b0; i7 = 1'b0; // testing 10000100    
    #50 i0 = 1'b0; i1 = 1'b1; i2 = 1'b1; i3 = 1'b1; i4 = 1'b1; i5 = 1'b1; i6 = 1'b1; i7 = 1'b1; // testing 01111111    
    
  end
  initial #950 $finish; //total time is 950 since 50 * 19 = 950 which is the total time needed for each input
endmodule
 
